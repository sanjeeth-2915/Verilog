module 4x1_mux ( input reg s0,s1,s2,a,b,c, output wire y);
  
