module sr_ff_tb;
  
