module 1:2_demux_tb;
reg sel;
  reg din;
  wire y0,y1;

  1:2
